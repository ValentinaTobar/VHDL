library verilog;
use verilog.vl_types.all;
entity ROM_128X8_SYNC_vlg_vec_tst is
end ROM_128X8_SYNC_vlg_vec_tst;
