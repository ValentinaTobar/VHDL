library verilog;
use verilog.vl_types.all;
entity output_ports_16_vlg_vec_tst is
end output_ports_16_vlg_vec_tst;
